module  y_ratio_case(data,raddr);
input        [10:0]     raddr;
output reg   [15:0]    data;

always@(*)
    case(raddr)
        11'd0   :   data  <=16'd40960;
        11'd1   :   data  <=16'hff99;
        11'd2   :   data  <=16'hff33;
        11'd3   :   data  <=16'hFECE;
        11'd4   :   data  <=16'hFE68;
        11'd5   :   data  <=16'hFE03;
        11'd6   :   data  <=16'hFD9F;
        11'd7   :   data  <=16'hFD3A;
        11'd8   :   data  <=16'hFCD6;
        11'd9   :   data  <=16'hFC73;
        11'd10   :   data <=16'hFC0F;

        11'd11   :   data <=16'hFBAC;
        11'd12   :   data <=16'hFB49;
        11'd13   :   data <=16'hFAE7;
        11'd14   :   data <=16'hFA85;
        11'd15   :   data <=16'hFA23;
        11'd16   :   data <=16'hF9C1;
        11'd17   :   data <=16'hF960;
        11'd18   :   data <=16'hF8FF;
        11'd19   :   data <=16'hF89E;
        11'd20   :   data <=16'hF83E;

        11'd21   :   data <=16'hF7DD;
        11'd22   :   data <=16'hF77E;
        11'd23   :   data <=16'hF71E;
        11'd24   :   data <=16'hF6BF;
        11'd25   :   data <=16'hF660;
        11'd26   :   data <=16'hF601;
        11'd27   :   data <=16'hF5A3;
        11'd28   :   data <=16'hF544;
        11'd29   :   data <=16'hF4E7;
        11'd30   :   data <=16'hF489;

        11'd31   :   data <=16'hF42C;
        11'd32   :   data <=16'hF3CF;
        11'd33   :   data <=16'hF372;
        11'd34   :   data <=16'hF316;
        11'd35   :   data <=16'hF2B9;
        11'd36   :   data <=16'hF25D;
        11'd37   :   data <=16'hF202;
        11'd38   :   data <=16'hF1A6;
        11'd39   :   data <=16'hF14B;
        11'd40   :   data <=16'hF0F0;

        11'd41   :   data <= 16'hF096;
        11'd42   :   data <= 16'hF03C;
        11'd43   :   data <= 16'hEFE2;
        11'd44   :   data <= 16'hEF88;
        11'd45   :   data <= 16'hEF2E;
        11'd46   :   data <= 16'hEED5;
        11'd47   :   data <= 16'hEE7C;
        11'd48   :   data <= 16'hEE23;
        11'd49   :   data <= 16'hEDCB;
        11'd50   :   data <= 16'hED73;

        11'd51   :   data <=16'hED1B;
        11'd52   :   data <=16'hECC3;
        11'd53   :   data <=16'hEC6B;
        11'd54   :   data <=16'hEC14;
        11'd55   :   data <=16'hEBBD;
        11'd56   :   data <=16'hEB66;
        11'd57   :   data <=16'hEB10;
        11'd58   :   data <=16'hEABA;
        11'd59   :   data <=16'hEA64;
        11'd60   :   data <=16'hEA0E;

        11'd61   :   data <=16'hE9B9;
        11'd62   :   data <=16'hE963;
        11'd63   :   data <=16'hE90E;
        11'd64   :   data <=16'hE8BA;
        11'd65   :   data <=16'hE865;
        11'd66   :   data <=16'hE811;
        11'd67   :   data <=16'hE7BD;
        11'd68   :   data <=16'hE769;
        11'd69   :   data <=16'hE716;
        11'd70   :   data <=16'hE6C2;

        11'd71   :   data <=16'hE66F;
        11'd72   :   data <=16'hE61C;
        11'd73   :   data <=16'hE5CA;
        11'd74   :   data <=16'hE577;
        11'd75   :   data <=16'hE525;
        11'd76   :   data <=16'hE4D3;
        11'd77   :   data <=16'hE481;
        11'd78   :   data <=16'hE430;
        11'd79   :   data <=16'hE3DF;
        11'd80   :   data <=16'hE38E;

        11'd81   :   data <=16'hE33D;
        11'd82   :   data <=16'hE2EC;
        11'd83   :   data <=16'hE29C;
        11'd84   :   data <=16'hE24C;
        11'd85   :   data <=16'hE1FC;
        11'd86   :   data <=16'hE1AC;
        11'd87   :   data <=16'hE15D;
        11'd88   :   data <=16'hE10E;
        11'd89   :   data <=16'hE0BF;
        11'd90   :   data <=16'hE070;

        11'd91   :   data <=16'hE021;
        11'd92   :   data <=16'hDFD3;
        11'd93   :   data <=16'hDF85;
        11'd94   :   data <=16'hDF37;
        11'd95   :   data <=16'hDEE9;
        11'd96   :   data <=16'hDE9B;
        11'd97   :   data <=16'hDE4E;
        11'd98   :   data <=16'hDE01;
        11'd99   :   data <=16'hDDB4;
        11'd100   :   data<=16'hDD67;

        11'd101   :   data <=16'hDD1B;
        11'd102   :   data <=16'hDCCF;
        11'd103   :   data <=16'hDC82;
        11'd104   :   data <=16'hDC37;
        11'd105   :   data <=16'hDBEB;
        11'd106   :   data <=16'hDB9F;
        11'd107   :   data <=16'hDB54;
        11'd108   :   data <=16'hDB09;
        11'd109   :   data <=16'hDABE;
        11'd110   :   data <=16'hDA74;

        11'd111   :   data <=16'hDA29;
        11'd112   :   data <=16'hD9DF;
        11'd113   :   data <=16'hD995;
        11'd114   :   data <=16'hD94B;
        11'd115   :   data <=16'hD901;
        11'd116   :   data <=16'hD8B8;
        11'd117   :   data <=16'hD86E;
        11'd118   :   data <=16'hD825;
        11'd119   :   data <=16'hD7DC;
        11'd120   :   data <=16'hD794;

        11'd121   :   data <=16'hD74B;
        11'd122   :   data <=16'hD703;
        11'd123   :   data <=16'hD6BB;
        11'd124   :   data <=16'hD673;
        11'd125   :   data <=16'hD62B;
        11'd126   :   data <=16'hD5E3;
        11'd127   :   data <=16'hD59C;
        11'd128   :   data <=16'hD555;
        11'd129   :   data <=16'hD50E;
        11'd130   :   data <=16'hD4C7;

        11'd131   :   data <=16'hD480;
        11'd132   :   data <=16'hD43A;
        11'd133   :   data <=16'hD3F4;
        11'd134   :   data <=16'hD3AD;
        11'd135   :   data <=16'hD368;
        11'd136   :   data <=16'hD322;
        11'd137   :   data <=16'hD2DC;
        11'd138   :   data <=16'hD297;
        11'd139   :   data <=16'hD252;
        11'd140   :   data <=16'hD20D;

        11'd141   :   data <=16'hD1C8;
        11'd142   :   data <=16'hD183;
        11'd143   :   data <=16'hD13F;
        11'd144   :   data <=16'hD0FA;
        11'd145   :   data <=16'hD0B6;
        11'd146   :   data <=16'hD072;
        11'd147   :   data <=16'hD02E;
        11'd148   :   data <=16'hCFEB;
        11'd149   :   data <=16'hCFA7;
        11'd150   :   data <=16'hCF64;

        11'd151   :   data <=16'hCF21;
        11'd152   :   data <=16'hCEDE;
        11'd153   :   data <=16'hCE9B;
        11'd154   :   data <=16'hCE58;
        11'd155   :   data <=16'hCE16;
        11'd156   :   data <=16'hCDD4;
        11'd157   :   data <=16'hCD92;
        11'd158   :   data <=16'hCD50;
        11'd159   :   data <=16'hCD0E;
        11'd160   :   data <=16'hCCCC;

        11'd161   :   data <=16'hCC8B;
        11'd162   :   data <=16'hCC4A;
        11'd163   :   data <=16'hCC08;
        11'd164   :   data <=16'hCBC7;
        11'd165   :   data <=16'hCB87;
        11'd166   :   data <=16'hCB46;
        11'd167   :   data <=16'hCB06;
        11'd168   :   data <=16'hCAC5;
        11'd169   :   data <=16'hCA85;
        11'd170   :   data <=16'hCA45;

        11'd171   :   data <=16'hCA05;
        11'd172   :   data <=16'hC9C5;
        11'd173   :   data <=16'hC986;
        11'd174   :   data <=16'hC947;
        11'd175   :   data <=16'hC907;
        11'd176   :   data <=16'hC8C8;
        11'd177   :   data <=16'hC889;
        11'd178   :   data <=16'hC84B;
        11'd179   :   data <=16'hC80C;
        11'd180   :   data <=16'hC7CE;

        11'd181   :   data <=16'hC78F;
        11'd182   :   data <=16'hC751;
        11'd183   :   data <=16'hC713;
        11'd184   :   data <=16'hC6D5;
        11'd185   :   data <=16'hC698;
        11'd186   :   data <=16'hC65A;
        11'd187   :   data <=16'hC61D;
        11'd188   :   data <=16'hC5DF;
        11'd189   :   data <=16'hC5A2;
        11'd190   :   data <=16'hC565;

        11'd191   :   data <=16'hC528;
        11'd192   :   data <=16'hC4EC;
        11'd193   :   data <=16'hC4AF;
        11'd194   :   data <=16'hC473;
        11'd195   :   data <=16'hC437;
        11'd196   :   data <=16'hC3FB;
        11'd197   :   data <=16'hC3BF;
        11'd198   :   data <=16'hC383;
        11'd199   :   data <=16'hC347;
        11'd200   :   data <=16'hC30C;

        11'd201   :   data <=16'hC2D0;
        11'd202   :   data <=16'hC295;
        11'd203   :   data <=16'hC25A;
        11'd204   :   data <=16'hC21F;
        11'd205   :   data <=16'hC1E4;
        11'd206   :   data <=16'hC1AA;
        11'd207   :   data <=16'hC16F;
        11'd208   :   data <=16'hC135;
        11'd209   :   data <=16'hC0FA;
        11'd210   :   data <=16'hC0C0;

        11'd211   :   data <=16'hC086;
        11'd212   :   data <=16'hC04C;
        11'd213   :   data <=16'hC013;
        11'd214   :   data <=16'hBFD9;
        11'd215   :   data <=16'hBFA0;
        11'd216   :   data <=16'hBF66;
        11'd217   :   data <=16'hBF2D;
        11'd218   :   data <=16'hBEF4;
        11'd219   :   data <=16'hBEBB;
        11'd220   :   data <=16'hBE82;

        11'd221   :   data <=16'hBE4A;
        11'd222   :   data <=16'hBE11;
        11'd223   :   data <=16'hBDD9;
        11'd224   :   data <=16'hBDA1;
        11'd225   :   data <=16'hBD69;
        11'd226   :   data <=16'hBD31;
        11'd227   :   data <=16'hBCF9;
        11'd228   :   data <=16'hBCC1;
        11'd229   :   data <=16'hBC89;
        11'd230   :   data <=16'hBC52;

        11'd231   :   data <=16'hBC1B;
        11'd232   :   data <=16'hBBE3;
        11'd233   :   data <=16'hBBAC;
        11'd234   :   data <=16'hBB75;
        11'd235   :   data <=16'hBB3E;
        11'd236   :   data <=16'hBB08;
        11'd237   :   data <=16'hBAD1;
        11'd238   :   data <=16'hBA9B;
        11'd239   :   data <=16'hBA64;
        11'd240   :   data <=16'hBA2E;

        11'd241   :   data <=16'hB9F8;
        11'd242   :   data <=16'hB9C2;
        11'd243   :   data <=16'hB98C;
        11'd244   :   data <=16'hB956;
        11'd245   :   data <=16'hB921;
        11'd246   :   data <=16'hB8EB;
        11'd247   :   data <=16'hB8B6;
        11'd248   :   data <=16'hB881;
        11'd249   :   data <=16'hB84C;
        11'd250   :   data <=16'hB817;


        11'd251   :   data <=16'hB7E2;
        11'd252   :   data <=16'hB7AD;
        11'd253   :   data <=16'hB778;
        11'd254   :   data <=16'hB744;
        11'd255   :   data <=16'hB70F;
        11'd256   :   data <=16'hB6DB;
        11'd257   :   data <=16'hB6A7;
        11'd258   :   data <=16'hB673;
        11'd259   :   data <=16'hB63F;
        11'd260   :   data <=16'hB60B;

        11'd261   :   data <=16'hB5D7;
        11'd262   :   data <=16'hB5A4;
        11'd263   :   data <=16'hB570;
        11'd264   :   data <=16'hB53D;
        11'd265   :   data <=16'hB509;
        11'd266   :   data <=16'hB4D6;
        11'd267   :   data <=16'hB4A3;
        11'd268   :   data <=16'hB470;
        11'd269   :   data <=16'hB43D;
        11'd270   :   data <=16'hB40B;

        11'd271   :   data <=16'hB3D8;
        11'd272   :   data <=16'hB3A6;
        11'd273   :   data <=16'hB373;
        11'd274   :   data <=16'hB341;
        11'd275   :   data <=16'hB30F;
        11'd276   :   data <=16'hB2DD;
        11'd277   :   data <=16'hB2AB;
        11'd278   :   data <=16'hB279;
        11'd279   :   data <=16'hB247;
        11'd280   :   data <=16'hB216;

        11'd281   :   data <=16'hB1E4;
        11'd282   :   data <=16'hB1B3;
        11'd283   :   data <=16'hB182;
        11'd284   :   data <=16'hB150;
        11'd285   :   data <=16'hB11F;
        11'd286   :   data <=16'hB0EE;
        11'd287   :   data <=16'hB0BD;
        11'd288   :   data <=16'hB08D;
        11'd289   :   data <=16'hB05C;
        11'd290   :   data <=16'hB02C;


        11'd291   :   data <=16'hAFFB;
        11'd292   :   data <=16'hAFCB;
        11'd293   :   data <=16'hAF9B;
        11'd294   :   data <=16'hAF6A;
        11'd295   :   data <=16'hAF3A;
        11'd296   :   data <=16'hAF0A;
        11'd297   :   data <=16'hAEDB;
        11'd298   :   data <=16'hAEAB;
        11'd299   :   data <=16'hAE7B;
        11'd300   :   data <=16'hAE4C;

        11'd301   :   data <=16'hAE1C;
        11'd302   :   data <=16'hADED;
        11'd303   :   data <=16'hADBE;
        11'd304   :   data <=16'hAD8F;
        11'd305   :   data <=16'hAD60;
        11'd306   :   data <=16'hAD31;
        11'd307   :   data <=16'hAD02;
        11'd308   :   data <=16'hACD3;
        11'd309   :   data <=16'hACA5;
        11'd310   :   data <=16'hAC76;

        11'd311   :   data <=16'hAC48;
        11'd312   :   data <=16'hAC19;
        11'd313   :   data <=16'hABEB;
        11'd314   :   data <=16'hABBD;
        11'd315   :   data <=16'hAB8F;
        11'd316   :   data <=16'hAB61;
        11'd317   :   data <=16'hAB33;
        11'd318   :   data <=16'hAB05;
        11'd319   :   data <=16'hAAD8;
        11'd320   :   data <=16'hAAAA;

        11'd321   :   data <=16'hAA7D;
        11'd322   :   data <=16'hAA4F;
        11'd323   :   data <=16'hAA22;
        11'd324   :   data <=16'hA9F5;
        11'd325   :   data <=16'hA9C8;
        11'd326   :   data <=16'hA99B;
        11'd327   :   data <=16'hA96E;
        11'd328   :   data <=16'hA941;
        11'd329   :   data <=16'hA914;
        11'd330   :   data <=16'hA8E8;

        11'd331   :   data <=16'hA8BB;
        11'd332   :   data <=16'hA88F;
        11'd333   :   data <=16'hA862;
        11'd334   :   data <=16'hA836;
        11'd335   :   data <=16'hA80A;
        11'd336   :   data <=16'hA7DE;
        11'd337   :   data <=16'hA7B2;
        11'd338   :   data <=16'hA786;
        11'd339   :   data <=16'hA75A;
        11'd340   :   data <=16'hA72F;

        11'd341   :   data <=16'hA703;
        11'd342   :   data <=16'hA6D7;
        11'd343   :   data <=16'hA6AC;
        11'd344   :   data <=16'hA681;
        11'd345   :   data <=16'hA655;
        11'd346   :   data <=16'hA62A;
        11'd347   :   data <=16'hA5FF;
        11'd348   :   data <=16'hA5D4;
        11'd349   :   data <=16'hA5A9;
        11'd350   :   data <=16'hA57E;

        11'd351   :   data <=16'hA553;
        11'd352   :   data <=16'hA529;
        11'd353   :   data <=16'hA4FE;
        11'd354   :   data <=16'hA4D4;
        11'd355   :   data <=16'hA4A9;
        11'd356   :   data <=16'hA47F;
        11'd357   :   data <=16'hA455;
        11'd358   :   data <=16'hA42B;
        11'd359   :   data <=16'hA401;
        11'd360   :   data <=16'hA3D7;

        11'd361   :   data <=16'hA3AD;
        11'd362   :   data <=16'hA383;
        11'd363   :   data <=16'hA359;
        11'd364   :   data <=16'hA32F;
        11'd365   :   data <=16'hA306;
        11'd366   :   data <=16'hA2DC;
        11'd367   :   data <=16'hA2B3;
        11'd368   :   data <=16'hA28A;
        11'd369   :   data <=16'hA260;
        11'd370   :   data <=16'hA237;

        11'd371   :   data <=16'hA20E;
        11'd372   :   data <=16'hA1E5;
        11'd373   :   data <=16'hA1BC;
        11'd374   :   data <=16'hA193;
        11'd375   :   data <=16'hA16B;
        11'd376   :   data <=16'hA142;
        11'd377   :   data <=16'hA119;
        11'd378   :   data <=16'hA0F1;
        11'd379   :   data <=16'hA0C8;
        11'd380   :   data <=16'hA0A0;

        11'd381   :   data <=16'hA078;
        11'd382   :   data <=16'hA050;
        11'd383   :   data <=16'hA028;
        11'd384   :   data <=16'hA000;
        11'd385   :   data <=16'h9FD8;
        11'd386   :   data <=16'h9FB0;
        11'd387   :   data <=16'h9F88;
        11'd388   :   data <=16'h9F60;
        11'd389   :   data <=16'h9F38;
        11'd390   :   data <=16'h9F11;

        11'd391   :   data <=16'h9EE9;
        11'd392   :   data <=16'h9EC2;
        11'd393   :   data <=16'h9E9B;
        11'd394   :   data <=16'h9E73;
        11'd395   :   data <=16'h9E4C;
        11'd396   :   data <=16'h9E25;
        11'd397   :   data <=16'h9DFE;
        11'd398   :   data <=16'h9DD7;
        11'd399   :   data <=16'h9DB0;
        11'd400   :   data <=16'h9D89;

        11'd401   :   data <=16'h9D63;
        11'd402   :   data <=16'h9D3C;
        11'd403   :   data <=16'h9D15;
        11'd404   :   data <=16'h9CEF;
        11'd405   :   data <=16'h9CC8;
        11'd406   :   data <=16'h9CA2;
        11'd407   :   data <=16'h9C7C;
        11'd408   :   data <=16'h9C55;
        11'd409   :   data <=16'h9C2F;
        11'd410   :   data <=16'h9C09;

        11'd411   :   data <=16'h9BE3;
        11'd412   :   data <=16'h9BBD;
        11'd413   :   data <=16'h9B97;
        11'd414   :   data <=16'h9B72;
        11'd415   :   data <=16'h9B4C;
        11'd416   :   data <=16'h9B26;
        11'd417   :   data <=16'h9B01;
        11'd418   :   data <=16'h9ADB;
        11'd419   :   data <=16'h9AB6;
        11'd420   :   data <=16'h9A90;

        11'd421   :   data <=16'h9A6B;
        11'd422   :   data <=16'h9A46;
        11'd423   :   data <=16'h9A21;
        11'd424   :   data <=16'h99FC;
        11'd425   :   data <=16'h99D7;
        11'd426   :   data <=16'h99B2;
        11'd427   :   data <=16'h998D;
        11'd428   :   data <=16'h9968;
        11'd429   :   data <=16'h9943;
        11'd430   :   data <=16'h991F;

        11'd431   :   data <=16'h98FA;
        11'd432   :   data <=16'h98D5;
        11'd433   :   data <=16'h98B1;
        11'd434   :   data <=16'h988D;
        11'd435   :   data <=16'h9868;
        11'd436   :   data <=16'h9844;
        11'd437   :   data <=16'h9820;
        11'd438   :   data <=16'h97FC;
        11'd439   :   data <=16'h97D8;
        11'd440   :   data <=16'h97B4;

        11'd441   :   data <=16'h9790;
        11'd442   :   data <=16'h976C;
        11'd443   :   data <=16'h9748;
        11'd444   :   data <=16'h9724;
        11'd445   :   data <=16'h9701;
        11'd446   :   data <=16'h96DD;
        11'd447   :   data <=16'h96BA;
        11'd448   :   data <=16'h9696;
        11'd449   :   data <=16'h9673;
        11'd450   :   data <=16'h964F;

        11'd451   :   data <=16'h962C;
        11'd452   :   data <=16'h9609;
        11'd453   :   data <=16'h95E6;
        11'd454   :   data <=16'h95C3;
        11'd455   :   data <=16'h95A0;
        11'd456   :   data <=16'h957D;
        11'd457   :   data <=16'h955A;
        11'd458   :   data <=16'h9537;
        11'd459   :   data <=16'h9514;
        11'd460   :   data <=16'h94F2;

        11'd461   :   data <=16'h94CF;
        11'd462   :   data <=16'h94AC;
        11'd463   :   data <=16'h948A;
        11'd464   :   data <=16'h9467;
        11'd465   :   data <=16'h9445;
        11'd466   :   data <=16'h9423;
        11'd467   :   data <=16'h9400;
        11'd468   :   data <=16'h93DE;
        11'd469   :   data <=16'h93BC;
        11'd470   :   data <=16'h939A;

        11'd471   :   data <=16'h9378;
        11'd472   :   data <=16'h9356;
        11'd473   :   data <=16'h9334;
        11'd474   :   data <=16'h9312;
        11'd475   :   data <=16'h92F1;
        11'd476   :   data <=16'h92CF;
        11'd477   :   data <=16'h92AD;
        11'd478   :   data <=16'h928C;
        11'd479   :   data <=16'h926A;
        11'd480   :   data <=16'h9249;

        11'd481   :   data <=16'h9227;
        11'd482   :   data <=16'h9206;
        11'd483   :   data <=16'h91E5;
        11'd484   :   data <=16'h91C3;
        11'd485   :   data <=16'h91A2;
        11'd486   :   data <=16'h9181;
        11'd487   :   data <=16'h9160;
        11'd488   :   data <=16'h913F;
        11'd489   :   data <=16'h911E;
        11'd490   :   data <=16'h90FD;

        11'd491   :   data <=16'h90DC;
        11'd492   :   data <=16'h90BC;
        11'd493   :   data <=16'h909B;
        11'd494   :   data <=16'h907A;
        11'd495   :   data <=16'h905A;
        11'd496   :   data <=16'h9039;
        11'd497   :   data <=16'h9019;
        11'd498   :   data <=16'h8FF8;
        11'd499   :   data <=16'h8FD8;
        11'd500   :   data <=16'h8FB8;

        11'd501   :   data <=16'h8F97;
        11'd502   :   data <=16'h8F77;
        11'd503   :   data <=16'h8F57;
        11'd504   :   data <=16'h8F37;
        11'd505   :   data <=16'h8F17;
        11'd506   :   data <=16'h8EF7;
        11'd507   :   data <=16'h8ED7;
        11'd508   :   data <=16'h8EB7;
        11'd509   :   data <=16'h8E97;
        11'd510   :   data <=16'h8E78;

        11'd511   :   data <=16'h8E58;
        11'd512   :   data <=16'h8E38;
        11'd513   :   data <=16'h8E19;
        11'd514   :   data <=16'h8DF9;
        11'd515   :   data <=16'h8DDA;
        11'd516   :   data <=16'h8DBA;
        11'd517   :   data <=16'h8D9B;
        11'd518   :   data <=16'h8D7C;
        11'd519   :   data <=16'h8D5C;
        11'd520   :   data <=16'h8D3D;

        11'd521   :   data <=16'h8D1E;
        11'd522   :   data <=16'h8CFF;
        11'd523   :   data <=16'h8CE0;
        11'd524   :   data <=16'h8CC1;
        11'd525   :   data <=16'h8CA2;
        11'd526   :   data <=16'h8C83;
        11'd527   :   data <=16'h8C64;
        11'd528   :   data <=16'h8C46;
        11'd529   :   data <=16'h8C27;
        11'd530   :   data <=16'h8C08;

        11'd531   :   data <=16'h8BEA;
        11'd532   :   data <=16'h8BCB;
        11'd533   :   data <=16'h8BAD;
        11'd534   :   data <=16'h8B8E;
        11'd535   :   data <=16'h8B70;
        11'd536   :   data <=16'h8B51;
        11'd537   :   data <=16'h8B33;
        11'd538   :   data <=16'h8B15;
        11'd539   :   data <=16'h8AF7;
        11'd540   :   data <=16'h8AD8;

        11'd541   :   data <=16'h8ABA;
        11'd542   :   data <=16'h8A9C;
        11'd543   :   data <=16'h8A7E;
        11'd544   :   data <=16'h8A60;
        11'd545   :   data <=16'h8A42;
        11'd546   :   data <=16'h8A25;
        11'd547   :   data <=16'h8A07;
        11'd548   :   data <=16'h89E9;
        11'd549   :   data <=16'h89CB;
        11'd550   :   data <=16'h89AE;

        11'd551   :   data <=16'h8990;
        11'd552   :   data <=16'h8973;
        11'd553   :   data <=16'h8955;
        11'd554   :   data <=16'h8938;
        11'd555   :   data <=16'h891A;
        11'd556   :   data <=16'h88FD;
        11'd557   :   data <=16'h88E0;
        11'd558   :   data <=16'h88C2;
        11'd559   :   data <=16'h88A5;
        11'd560   :   data <=16'h8888;

        11'd561   :   data <=16'h886B;
        11'd562   :   data <=16'h884E;
        11'd563   :   data <=16'h8831;
        11'd564   :   data <=16'h8814;
        11'd565   :   data <=16'h87F7;
        11'd566   :   data <=16'h87DA;
        11'd567   :   data <=16'h87BD;
        11'd568   :   data <=16'h87A1;
        11'd569   :   data <=16'h8784;
        11'd570   :   data <=16'h8767;

        11'd571   :   data <=16'h874B;
        11'd572   :   data <=16'h872E;
        11'd573   :   data <=16'h8711;
        11'd574   :   data <=16'h86F5;
        11'd575   :   data <=16'h86D9;
        11'd576   :   data <=16'h86BC;
        11'd577   :   data <=16'h86A0;
        11'd578   :   data <=16'h8683;
        11'd579   :   data <=16'h8667;
        11'd580   :   data <=16'h864B;

        11'd581   :   data <=16'h862F;
        11'd582   :   data <=16'h8613;
        11'd583   :   data <=16'h85F7;
        11'd584   :   data <=16'h85DB;
        11'd585   :   data <=16'h85BF;
        11'd586   :   data <=16'h85A3;
        11'd587   :   data <=16'h8587;
        11'd588   :   data <=16'h856B;
        11'd589   :   data <=16'h854F;
        11'd590   :   data <=16'h8534;

        11'd591   :   data <=16'h8518;
        11'd592   :   data <=16'h84FC;
        11'd593   :   data <=16'h84E1;
        11'd594   :   data <=16'h84C5;
        11'd595   :   data <=16'h84A9;
        11'd596   :   data <=16'h848E;
        11'd597   :   data <=16'h8473;
        11'd598   :   data <=16'h8457;
        11'd599   :   data <=16'h843C;
        11'd600   :   data <=16'h8421;

        11'd601   :   data <=16'h8405;
        11'd602   :   data <=16'h83EA;
        11'd603   :   data <=16'h83CF;
        11'd604   :   data <=16'h83B4;
        11'd605   :   data <=16'h8399;
        11'd606   :   data <=16'h837E;
        11'd607   :   data <=16'h8363;
        11'd608   :   data <=16'h8348;
        11'd609   :   data <=16'h832D;
        11'd610   :   data <=16'h8312;

        11'd611   :   data <=16'h82F7;
        11'd612   :   data <=16'h82DC;
        11'd613   :   data <=16'h82C2;
        11'd614   :   data <=16'h82A7;
        11'd615   :   data <=16'h828C;
        11'd616   :   data <=16'h8272;
        11'd617   :   data <=16'h8257;
        11'd618   :   data <=16'h823D;
        11'd619   :   data <=16'h8222;
        11'd620   :   data <=16'h8208;

        11'd621   :   data <=16'h81ED;
        11'd622   :   data <=16'h81D3;
        11'd623   :   data <=16'h81B9;
        11'd624   :   data <=16'h819E;
        11'd625   :   data <=16'h8184;
        11'd626   :   data <=16'h816A;
        11'd627   :   data <=16'h8150;
        11'd628   :   data <=16'h8136;
        11'd629   :   data <=16'h811C;
        11'd630   :   data <=16'h8102;

        11'd631   :   data <=16'h80E8;
        11'd632   :   data <=16'h80CE;
        11'd633   :   data <=16'h80B4;
        11'd634   :   data <=16'h809A;
        11'd635   :   data <=16'h8080;
        11'd636   :   data <=16'h8066;
        11'd637   :   data <=16'h804C;
        11'd638   :   data <=16'h8033;
        11'd639   :   data <=16'h8019;
        11'd640  :   data <= 16'h8000;

        11'd641   :   data <=16'h7FE6;
        11'd642   :   data <=16'h7FCC;
        11'd643   :   data <=16'h7FB3;
        11'd644   :   data <=16'h7F99;
        11'd645   :   data <=16'h7F80;
        11'd646   :   data <=16'h7F67;
        11'd647   :   data <=16'h7F4D;
        11'd648   :   data <=16'h7F34;
        11'd649   :   data <=16'h7F1B;
        11'd650  :   data <= 16'h7F01;

        11'd651   :   data <=16'h7EE8;
        11'd652   :   data <=16'h7ECF;
        11'd653   :   data <=16'h7EB6;
        11'd654   :   data <=16'h7E9D;
        11'd655   :   data <=16'h7E84;
        11'd656   :   data <=16'h7E6B;
        11'd657   :   data <=16'h7E52;
        11'd658   :   data <=16'h7E39;
        11'd659   :   data <=16'h7E20;
        11'd660  :   data <= 16'h7E07;

        11'd661   :   data <=16'h7DEF;
        11'd662   :   data <=16'h7DD6;
        11'd663   :   data <=16'h7DBD;
        11'd664   :   data <=16'h7DA4;
        11'd665   :   data <=16'h7D8C;
        11'd666   :   data <=16'h7D73;
        11'd667   :   data <=16'h7D5B;
        11'd668   :   data <=16'h7D42;
        11'd669   :   data <=16'h7D2A;
        11'd670  :   data <= 16'h7D11;

        11'd671   :   data <=16'h7CF9;
        11'd672   :   data <=16'h7CE0;
        11'd673   :   data <=16'h7CC8;
        11'd674   :   data <=16'h7CB0;
        11'd675   :   data <=16'h7C97;
        11'd676   :   data <=16'h7C7F;
        11'd677   :   data <=16'h7C67;
        11'd678   :   data <=16'h7C4F;
        11'd679   :   data <=16'h7C37;
        11'd680  :   data <= 16'h7C1F;

        11'd681   :   data <=16'h7C06;
        11'd682   :   data <=16'h7BEE;
        11'd683   :   data <=16'h7BD6;
        11'd684   :   data <=16'h7BBF;
        11'd685   :   data <=16'h7BA7;
        11'd686   :   data <=16'h7B8F;
        11'd687   :   data <=16'h7B77;
        11'd688   :   data <=16'h7B5F;
        11'd689   :   data <=16'h7B47;
        11'd690  :   data <= 16'h7B30;

        11'd691   :   data <=16'h7B18;
        11'd692   :   data <=16'h7B00;
        11'd693   :   data <=16'h7AE9;
        11'd694   :   data <=16'h7AD1;
        11'd695   :   data <=16'h7ABA;
        11'd696   :   data <=16'h7AA2;
        11'd697   :   data <=16'h7A8B;
        11'd698   :   data <=16'h7A73;
        11'd699   :   data <=16'h7A5C;
        11'd700  :   data <= 16'h7A44;

        11'd701   :   data <=16'h7A2D;
        11'd702   :   data <=16'h7A16;
        11'd703   :   data <=16'h79FE;
        11'd704   :   data <=16'h79E7;
        11'd705   :   data <=16'h79D0;
        11'd706   :   data <=16'h79B9;
        11'd707   :   data <=16'h79A2;
        11'd708   :   data <=16'h798B;
        11'd709   :   data <=16'h7973;
        11'd710  :   data <= 16'h795C;

        11'd711   :   data <=16'h7945;
        11'd712   :   data <=16'h792E;
        11'd713   :   data <=16'h7918;
        11'd714   :   data <=16'h7901;
        11'd715   :   data <=16'h78EA;
        11'd716   :   data <=16'h78D3;
        11'd717   :   data <=16'h78BC;
        11'd718   :   data <=16'h78A5;
        11'd719   :   data <=16'h788F;
        11'd720  :   data <= 16'h7878;

        11'd721   :   data <=16'h7861;
        11'd722   :   data <=16'h784B;
        11'd723   :   data <=16'h7834;
        11'd724   :   data <=16'h781E;
        11'd725   :   data <=16'h7807;
        11'd726   :   data <=16'h77F1;
        11'd727   :   data <=16'h77DA;
        11'd728   :   data <=16'h77C4;
        11'd729   :   data <=16'h77AD;
        11'd730  :   data <= 16'h7797;

        11'd731   :   data <=16'h7781;
        11'd732   :   data <=16'h776A;
        11'd733   :   data <=16'h7754;
        11'd734   :   data <=16'h773E;
        11'd735   :   data <=16'h7728;
        11'd736   :   data <=16'h7711;
        11'd737   :   data <=16'h76FB;
        11'd738   :   data <=16'h76E5;
        11'd739   :   data <=16'h76CF;
        11'd740  :   data <= 16'h76B9;

        11'd741   :   data <=16'h76A3;
        11'd742   :   data <=16'h768D;
        11'd743   :   data <=16'h7677;
        11'd744   :   data <=16'h7661;
        11'd745   :   data <=16'h764B;
        11'd746   :   data <=16'h7635;
        11'd747   :   data <=16'h7620;
        11'd748   :   data <=16'h760A;
        11'd749   :   data <=16'h75F4;
        11'd750  :   data <= 16'h75DE;

        11'd751   :   data <=16'h75C9;
        11'd752   :   data <=16'h75B3;
        11'd753   :   data <=16'h759D;
        11'd754   :   data <=16'h7588;
        11'd755   :   data <=16'h7572;
        11'd756   :   data <=16'h755D;
        11'd757   :   data <=16'h7547;
        11'd758   :   data <=16'h7532;
        11'd759   :   data <=16'h751C;
        11'd760  :   data <= 16'h7507;

        11'd761   :   data <=16'h74F1;
        11'd762   :   data <=16'h74DC;
        11'd763   :   data <=16'h74C7;
        11'd764   :   data <=16'h74B1;
        11'd765   :   data <=16'h749C;
        11'd766   :   data <=16'h7487;
        11'd767   :   data <=16'h7472;
        11'd768   :   data <=16'h745D;
        11'd769   :   data <=16'h7447;
        11'd770  :   data <= 16'h7432;

        11'd771   :   data <=16'h741D;
        11'd772   :   data <=16'h7408;
        11'd773   :   data <=16'h73F3;
        11'd774   :   data <=16'h73DE;
        11'd775   :   data <=16'h73C9;
        11'd776   :   data <=16'h73B4;
        11'd777   :   data <=16'h739F;
        11'd778   :   data <=16'h738B;
        11'd779   :   data <=16'h7376;
        11'd780  :   data <= 16'h7361;

        11'd781   :   data <=16'h734C;
        11'd782   :   data <=16'h7337;
        11'd783   :   data <=16'h7323;
        11'd784   :   data <=16'h730E;
        11'd785   :   data <=16'h72F9;
        11'd786   :   data <=16'h72E5;
        11'd787   :   data <=16'h72D0;
        11'd788   :   data <=16'h72BB;
        11'd789   :   data <=16'h72A7;
        11'd790  :   data <= 16'h7292;

        11'd791   :   data <=16'h80E8;
        11'd792   :   data <=16'h80CE;
        11'd793   :   data <=16'h80B4;
        11'd794   :   data <=16'h809A;
        11'd795   :   data <=16'h8080;
        11'd796   :   data <=16'h8066;
        11'd797   :   data <=16'h804C;
        11'd798   :   data <=16'h8033;
        11'd799   :   data <=16'h8019;
        11'd800  :   data <= 16'h8000;

        11'd801   :   data <=16'h71B2;
        11'd802   :   data <=16'h719E;
        11'd803   :   data <=16'h718A;
        11'd804   :   data <=16'h7176;
        11'd805   :   data <=16'h7162;
        11'd806   :   data <=16'h714E;
        11'd807   :   data <=16'h713A;
        11'd808   :   data <=16'h7126;
        11'd809   :   data <=16'h7112;
        11'd810   :   data <=16'h70FE;

        11'd811   :   data <=16'h70EA;
        11'd812   :   data <=16'h70D6;
        11'd813   :   data <=16'h70C2;
        11'd814   :   data <=16'h70AE;
        11'd815   :   data <=16'h709A;
        11'd816   :   data <=16'h7087;
        11'd817   :   data <=16'h7073;
        11'd818   :   data <=16'h705F;
        11'd819   :   data <=16'h704B;
        11'd820   :   data <=16'h7038;

        11'd821   :   data <=16'h7024;
        11'd822   :   data <=16'h7010;
        11'd823   :   data <=16'h6FFD;
        11'd824   :   data <=16'h6FE9;
        11'd825   :   data <=16'h6FD6;
        11'd826   :   data <=16'h6FC2;
        11'd827   :   data <=16'h6FAF;
        11'd828   :   data <=16'h6F9B;
        11'd829   :   data <=16'h6F88;
        11'd830   :   data <=16'h6F74;

        11'd831   :   data <=16'h6F61;
        11'd832   :   data <=16'h6F4D;
        11'd833   :   data <=16'h6F3A;
        11'd834   :   data <=16'h6F27;
        11'd835   :   data <=16'h6F13;
        11'd836   :   data <=16'h6F00;
        11'd837   :   data <=16'h6EED;
        11'd838   :   data <=16'h6EDA;
        11'd839   :   data <=16'h6EC7;
        11'd840   :   data <=16'h6EB3;

        11'd841   :   data <=16'h6EA0;
        11'd842   :   data <=16'h6E8D;
        11'd843   :   data <=16'h6E7A;
        11'd844   :   data <=16'h6E67;
        11'd845   :   data <=16'h6E54;
        11'd846   :   data <=16'h6E41;
        11'd847   :   data <=16'h6E2E;
        11'd848   :   data <=16'h6E1B;
        11'd849   :   data <=16'h6E08;
        11'd850   :   data <=16'h6DF5;

        11'd851   :   data <=16'h6DE2;
        11'd852   :   data <=16'h6DCF;
        11'd853   :   data <=16'h6DBD;
        11'd854   :   data <=16'h6DAA;
        11'd855   :   data <=16'h6D97;
        11'd856   :   data <=16'h6D84;
        11'd857   :   data <=16'h6D72;
        11'd858   :   data <=16'h6D5F;
        11'd859   :   data <=16'h6D4C;
        11'd860   :   data <=16'h6D3A;

        11'd861   :   data <=16'h6D27;
        11'd862   :   data <=16'h6D14;
        11'd863   :   data <=16'h6D02;
        11'd864   :   data <=16'h6CEF;
        11'd865   :   data <=16'h6CDD;
        11'd866   :   data <=16'h6CCA;
        11'd867   :   data <=16'h6CB8;
        11'd868   :   data <=16'h6CA5;
        11'd869   :   data <=16'h6C93;
        11'd870   :   data <=16'h6C80;

        11'd871   :   data <=16'h6C6E;
        11'd872   :   data <=16'h6C5C;
        11'd873   :   data <=16'h6C49;
        11'd874   :   data <=16'h6C37;
        11'd875   :   data <=16'h6C25;
        11'd876   :   data <=16'h6C12;
        11'd877   :   data <=16'h6C00;
        11'd878   :   data <=16'h6BEE;
        11'd879   :   data <=16'h6BDC;
        11'd880   :   data <=16'h6BCA;

        11'd881   :   data <=16'h6BB7;
        11'd882   :   data <=16'h6BA5;
        11'd883   :   data <=16'h6B93;
        11'd884   :   data <=16'h6B81;
        11'd885   :   data <=16'h6B6F;
        11'd886   :   data <=16'h6B5D;
        11'd887   :   data <=16'h6B4B;
        11'd888   :   data <=16'h6B39;
        11'd889   :   data <=16'h6B27;
        11'd890   :   data <=16'h6B15;

        11'd891   :   data <=16'h6B03;
        11'd892   :   data <=16'h6AF1;
        11'd893   :   data <=16'h6AE0;
        11'd894   :   data <=16'h6ACE;
        11'd895   :   data <=16'h6ABC;
        11'd896   :   data <=16'h6AAA;
        11'd897   :   data <=16'h6A98;
        11'd898   :   data <=16'h6A87;
        11'd899   :   data <=16'h6A75;
        11'd900   :   data <=16'h6A63;

        11'd901   :   data <=16'h6A52;
        11'd902   :   data <=16'h6A40;
        11'd903   :   data <=16'h6A2E;
        11'd904   :   data <=16'h6A1D;
        11'd905   :   data <=16'h6A0B;
        11'd906   :   data <=16'h69FA;
        11'd907   :   data <=16'h69E8;
        11'd908   :   data <=16'h69D6;
        11'd909   :   data <=16'h69C5;
        11'd910   :   data <=16'h69B4;

        11'd911   :   data <=16'h69A2;
        11'd912   :   data <=16'h6991;
        11'd913   :   data <=16'h697F;
        11'd914   :   data <=16'h696E;
        11'd915   :   data <=16'h695D;
        11'd916   :   data <=16'h694B;
        11'd917   :   data <=16'h693A;
        11'd918   :   data <=16'h6929;
        11'd919   :   data <=16'h6917;
        11'd920   :   data <=16'h6906;

        11'd921   :   data <=16'h68F5;
        11'd922   :   data <=16'h68E4;
        11'd923   :   data <=16'h68D2;
        11'd924   :   data <=16'h68C1;
        11'd925   :   data <=16'h68B0;
        11'd926   :   data <=16'h689F;
        11'd927   :   data <=16'h688E;
        11'd928   :   data <=16'h687D;
        11'd929   :   data <=16'h686C;
        11'd930   :   data <=16'h685B;

        11'd921   :   data <=16'h68F5;
        11'd922   :   data <=16'h68E4;
        11'd923   :   data <=16'h68D2;
        11'd924   :   data <=16'h68C1;
        11'd925   :   data <=16'h68B0;
        11'd926   :   data <=16'h689F;
        11'd927   :   data <=16'h688E;
        11'd928   :   data <=16'h687D;
        11'd929   :   data <=16'h686C;
        11'd930   :   data <=16'h685B;

        11'd931   :   data <=16'h684A;
        11'd932   :   data <=16'h6839;
        11'd933   :   data <=16'h6828;
        11'd934   :   data <=16'h6817;
        11'd935   :   data <=16'h6806;
        11'd936   :   data <=16'h67F5;
        11'd937   :   data <=16'h67E4;
        11'd938   :   data <=16'h67D3;
        11'd939   :   data <=16'h67C3;
        11'd940   :   data <=16'h67B2;

        11'd941   :   data <=16'h67A1;
        11'd942   :   data <=16'h6790;
        11'd943   :   data <=16'h677F;
        11'd944   :   data <=16'h676F;
        11'd945   :   data <=16'h675E;
        11'd946   :   data <=16'h674D;
        11'd947   :   data <=16'h673D;
        11'd948   :   data <=16'h672C;
        11'd949   :   data <=16'h671B;
        11'd950   :   data <=16'h670B;

        11'd951   :   data <=16'h66FA;
        11'd952   :   data <=16'h66EA;
        11'd953   :   data <=16'h66D9;
        11'd954   :   data <=16'h66C9;
        11'd955   :   data <=16'h66B8;
        11'd956   :   data <=16'h66A8;
        11'd957   :   data <=16'h6697;
        11'd958   :   data <=16'h6687;
        11'd959   :   data <=16'h6676;
        11'd960   :   data <=16'h6666;

        11'd961   :   data <=16'h6656;
        11'd962   :   data <=16'h6645;
        11'd963   :   data <=16'h6635;
        11'd964   :   data <=16'h6625;
        11'd965   :   data <=16'h6614;
        11'd966   :   data <=16'h6604;
        11'd967   :   data <=16'h65F4;
        11'd968   :   data <=16'h65E3;
        11'd969   :   data <=16'h65D3;
        11'd970   :   data <=16'h65C3;

        11'd971   :   data <=16'h65B3;
        11'd972   :   data <=16'h65A3;
        11'd973   :   data <=16'h6593;
        11'd974   :   data <=16'h6583;
        11'd975   :   data <=16'h6572;
        11'd976   :   data <=16'h6562;
        11'd977   :   data <=16'h6552;
        11'd978   :   data <=16'h6542;
        11'd979   :   data <=16'h6532;
        11'd980   :   data <=16'h6522;

        11'd981   :   data <=16'h6512;
        11'd982   :   data <=16'h6502;
        11'd983   :   data <=16'h64F2;
        11'd984   :   data <=16'h64E2;
        11'd985   :   data <=16'h64D3;
        11'd986   :   data <=16'h64C3;
        11'd987   :   data <=16'h64B3;
        11'd988   :   data <=16'h64A3;
        11'd989   :   data <=16'h6493;
        11'd990   :   data <=16'h6483;

        11'd991   :   data <=16'h6474;
        11'd992   :   data <=16'h6464;
        11'd993   :   data <=16'h6454;
        11'd994   :   data <=16'h6444;
        11'd995   :   data <=16'h6435;
        11'd996   :   data <=16'h6425;
        11'd997   :   data <=16'h6415;
        11'd998   :   data <=16'h6406;
        11'd999   :   data <=16'h63F6;
        11'd1000  :   data <=16'h63E7;

        11'd1001   :   data  <=16'h63D7;
        11'd1002   :   data  <=16'h63C7;
        11'd1003   :   data  <=16'h63B8;
        11'd1004   :   data  <=16'h63A8;
        11'd1005   :   data  <=16'h6399;
        11'd1006   :   data  <=16'h6389;
        11'd1007   :   data  <=16'h637A;
        11'd1008   :   data  <=16'h636A;
        11'd1009   :   data  <=16'h635B;
        11'd1010   :   data  <=16'h634C;

        11'd1011   :   data <=16'h633C;
        11'd1012   :   data <=16'h632D;
        11'd1013   :   data <=16'h631D;
        11'd1014   :   data <=16'h630E;
        11'd1015   :   data <=16'h62FF;
        11'd1016   :   data <=16'h62EF;
        11'd1017   :   data <=16'h62E0;
        11'd1018   :   data <=16'h62D1;
        11'd1019   :   data <=16'h62C2;
        11'd1020   :   data <=16'h62B2;

        11'd1021   :   data <=16'h62A3;
        11'd1022   :   data <=16'h6294;
        11'd1023   :   data <=16'h6285;
        11'd1024   :   data <=16'h6276;
        11'd1025   :   data <=16'h6267;
        11'd1026   :   data <=16'h6257;
        11'd1027   :   data <=16'h6248;
        11'd1028   :   data <=16'h6239;
        11'd1029   :   data <=16'h622A;
        11'd1030   :   data <=16'h621B;

        11'd1031   :   data <=16'h620C;
        11'd1032   :   data <=16'h61FD;
        11'd1033   :   data <=16'h61EE;
        11'd1034   :   data <=16'h61DF;
        11'd1035   :   data <=16'h61D0;
        11'd1036   :   data <=16'h61C1;
        11'd1037   :   data <=16'h61B2;
        11'd1038   :   data <=16'h61A3;
        11'd1039   :   data <=16'h6194;
        11'd1040   :   data <=16'h6186;

        11'd1041   :   data <= 16'h6177;
        11'd1042   :   data <= 16'h6168;
        11'd1043   :   data <= 16'h6159;
        11'd1044   :   data <= 16'h614A;
        11'd1045   :   data <= 16'h613C;
        11'd1046   :   data <= 16'h612D;
        11'd1047   :   data <= 16'h611E;
        11'd1048   :   data <= 16'h610F;
        11'd1049   :   data <= 16'h6101;
        11'd1050   :   data <= 16'h60F2;

        11'd1051   :   data <=16'h60E3;
        11'd1052   :   data <=16'h60D5;
        11'd1053   :   data <=16'h60C6;
        11'd1054   :   data <=16'h60B7;
        11'd1055   :   data <=16'h60A9;
        11'd1056   :   data <=16'h609A;
        11'd1057   :   data <=16'h608B;
        11'd1058   :   data <=16'h607D;
        11'd1059   :   data <=16'h606E;
        11'd1060   :   data <=16'h6060;

        11'd1061   :   data <=16'h6051;
        11'd1062   :   data <=16'h6043;
        11'd1063   :   data <=16'h6034;
        11'd1064   :   data <=16'h6026;
        11'd1065   :   data <=16'h6018;
        11'd1066   :   data <=16'h6009;
        11'd1067   :   data <=16'h5FFB;
        11'd1068   :   data <=16'h5FEC;
        11'd1069   :   data <=16'h5FDE;
        11'd1070   :   data <=16'h5FD0;

        11'd1071   :   data <=16'h5FC1;
        11'd1072   :   data <=16'h5FB3;
        11'd1073   :   data <=16'h5FA5;
        11'd1074   :   data <=16'h5F96;
        11'd1075   :   data <=16'h5F88;
        11'd1076   :   data <=16'h5F7A;
        11'd1077   :   data <=16'h5F6C;
        11'd1078   :   data <=16'h5F5D;
        11'd1079   :   data <=16'h5F4F;
        11'd1080   :   data <=16'h5F41;

        11'd1081   :   data <=16'h5F33;
        11'd1082   :   data <=16'h5F25;
        11'd1083   :   data <=16'h5F17;
        11'd1084   :   data <=16'h5F08;
        11'd1085   :   data <=16'h5EFA;
        11'd1086   :   data <=16'h5EEC;
        11'd1087   :   data <=16'h5EDE;
        11'd1088   :   data <=16'h5ED0;
        11'd1089   :   data <=16'h5EC2;
        11'd1090   :   data <=16'h5EB4;

        11'd1091   :   data <=16'h5EA6;
        11'd1092   :   data <=16'h5E98;
        11'd1093   :   data <=16'h5E8A;
        11'd1094   :   data <=16'h5E7C;
        11'd1095   :   data <=16'h5E6E;
        11'd1096   :   data <=16'h5E60;
        11'd1097   :   data <=16'h5E52;
        11'd1098   :   data <=16'h5E44;
        11'd1099   :   data <=16'h5E37;
        11'd1100   :   data<= 16'h5E29;

        11'd1101   :   data  <=16'h5E1B;
        11'd1102   :   data  <=16'h5E0D;
        11'd1103   :   data  <=16'h5DFF;
        11'd1104   :   data  <=16'h5DF1;
        11'd1105   :   data  <=16'h5DE4;
        11'd1106   :   data  <=16'h5DD6;
        11'd1107   :   data  <=16'h5DC8;
        11'd1108   :   data  <=16'h5DBA;
        11'd1109   :   data  <=16'h5DAD;
        11'd1110   :   data  <=16'h5D9F;

        11'd1111   :   data <=16'h5D91;
        11'd1112   :   data <=16'h5D84;
        11'd1113   :   data <=16'h5D76;
        11'd1114   :   data <=16'h5D68;
        11'd1115   :   data <=16'h5D5B;
        11'd1116   :   data <=16'h5D4D;
        11'd1117   :   data <=16'h5D3F;
        11'd1118   :   data <=16'h5D32;
        11'd1119   :   data <=16'h5D24;
        11'd1120   :   data <=16'h5D17;

        11'd1121   :   data <=16'h5D09;
        11'd1122   :   data <=16'h5CFC;
        11'd1123   :   data <=16'h5CEE;
        11'd1124   :   data <=16'h5CE1;
        11'd1125   :   data <=16'h5CD3;
        11'd1126   :   data <=16'h5CC6;
        11'd1127   :   data <=16'h5CB8;
        11'd1128   :   data <=16'h5CAB;
        11'd1129   :   data <=16'h5C9E;
        11'd1130   :   data <=16'h5C90;

        11'd1131   :   data <=16'h5C83;
        11'd1132   :   data <=16'h5C75;
        11'd1133   :   data <=16'h5C68;
        11'd1134   :   data <=16'h5C5B;
        11'd1135   :   data <=16'h5C4D;
        11'd1136   :   data <=16'h5C40;
        11'd1137   :   data <=16'h5C33;
        11'd1138   :   data <=16'h5C26;
        11'd1139   :   data <=16'h5C18;
        11'd1140   :   data <=16'h5C0B;

        11'd1141   :   data <= 16'h5BFE;
        11'd1142   :   data <= 16'h5BF1;
        11'd1143   :   data <= 16'h5BE3;
        11'd1144   :   data <= 16'h5BD6;
        11'd1145   :   data <= 16'h5BC9;
        11'd1146   :   data <= 16'h5BBC;
        11'd1147   :   data <= 16'h5BAF;
        11'd1148   :   data <= 16'h5BA2;
        11'd1149   :   data <= 16'h5B94;
        11'd1150   :   data <= 16'h5B87;

        11'd1151   :   data <=16'hED1B;
        11'd1152   :   data <=16'hECC3;
        11'd1153   :   data <=16'hEC6B;
        11'd1154   :   data <=16'hEC14;
        11'd1155   :   data <=16'hEBBD;
        11'd1156   :   data <=16'hEB66;
        11'd1157   :   data <=16'hEB10;
        11'd1158   :   data <=16'hEABA;
        11'd1159   :   data <=16'hEA64;
        11'd1160   :   data <=16'hEA0E;

        11'd1161   :   data <=16'h5AF8;
        11'd1162   :   data <=16'h5AEB;
        11'd1163   :   data <=16'h5ADE;
        11'd1164   :   data <=16'h5AD2;
        11'd1165   :   data <=16'h5AC5;
        11'd1166   :   data <=16'h5AB8;
        11'd1167   :   data <=16'h5AAB;
        11'd1168   :   data <=16'h5A9E;
        11'd1169   :   data <=16'h5A91;
        11'd1170   :   data <=16'h5A84;

        11'd1171   :   data <=16'h5A78;
        11'd1172   :   data <=16'h5A6B;
        11'd1173   :   data <=16'h5A5E;
        11'd1174   :   data <=16'h5A51;
        11'd1175   :   data <=16'h5A45;
        11'd1176   :   data <=16'h5A38;
        11'd1177   :   data <=16'h5A2B;
        11'd1178   :   data <=16'h5A1E;
        11'd1179   :   data <=16'h5A12;
        11'd1180   :   data <=16'h5A05;

        11'd1181   :   data <=16'h59F8;
        11'd1182   :   data <=16'h59EC;
        11'd1183   :   data <=16'h59DF;
        11'd1184   :   data <=16'h59D3;
        11'd1185   :   data <=16'h59C6;
        11'd1186   :   data <=16'h59B9;
        11'd1187   :   data <=16'h59AD;
        11'd1188   :   data <=16'h59A0;
        11'd1189   :   data <=16'h5994;
        11'd1190   :   data <=16'h5987;

        11'd1191   :   data <=16'h597B;
        11'd1192   :   data <=16'h596E;
        11'd1193   :   data <=16'h5962;
        11'd1194   :   data <=16'h5955;
        11'd1195   :   data <=16'h5949;
        11'd1196   :   data <=16'h593C;
        11'd1197   :   data <=16'h5930;
        11'd1198   :   data <=16'h5923;
        11'd1199   :   data <=16'h5917;
        11'd1200   :   data<= 16'h590B;

        11'd1201   :   data  <=16'h58FE;
        11'd1202   :   data  <=16'h58F2;
        11'd1203   :   data  <=16'h58E6;
        11'd1204   :   data  <=16'h58D9;
        11'd1205   :   data  <=16'h58CD;
        11'd1206   :   data  <=16'h58C1;
        11'd1207   :   data  <=16'h58B4;
        11'd1208   :   data  <=16'h58A8;
        11'd1209   :   data  <=16'h589C;
        11'd1210   :   data  <=16'h588F;

        11'd1211   :   data <=16'h5883;
        11'd1212   :   data <=16'h5877;
        11'd1213   :   data <=16'h586B;
        11'd1214   :   data <=16'h585E;
        11'd1215   :   data <=16'h5852;
        11'd1216   :   data <=16'h5846;
        11'd1217   :   data <=16'h583A;
        11'd1218   :   data <=16'h582E;
        11'd1219   :   data <=16'h5822;
        11'd1220   :   data <=16'h5816;

        11'd1221   :   data <=16'h5809;
        11'd1222   :   data <=16'h57FD;
        11'd1223   :   data <=16'h57F1;
        11'd1224   :   data <=16'h57E5;
        11'd1225   :   data <=16'h57D9;
        11'd1226   :   data <=16'h57CD;
        11'd1227   :   data <=16'h57C1;
        11'd1228   :   data <=16'h57B5;
        11'd1229   :   data <=16'h57A9;
        11'd1230   :   data <=16'h579D;

        11'd1231   :   data <=16'h5791;
        11'd1232   :   data <=16'h5785;
        11'd1233   :   data <=16'h5779;
        11'd1234   :   data <=16'h576D;
        11'd1235   :   data <=16'h5761;
        11'd1236   :   data <=16'h5755;
        11'd1237   :   data <=16'h5749;
        11'd1238   :   data <=16'h573D;
        11'd1239   :   data <=16'h5732;
        11'd1240   :   data <=16'h5726;

        11'd1241   :   data <= 16'h571A;
        11'd1242   :   data <= 16'h570E;
        11'd1243   :   data <= 16'h5702;
        11'd1244   :   data <= 16'h56F6;
        11'd1245   :   data <= 16'h56EA;
        11'd1246   :   data <= 16'h56DF;
        11'd1247   :   data <= 16'h56D3;
        11'd1248   :   data <= 16'h56C7;
        11'd1249   :   data <= 16'h56BB;
        11'd1250   :   data <= 16'h56B0;

        11'd1251   :   data <=16'h56A4;
        11'd1252   :   data <=16'h5698;
        11'd1253   :   data <=16'h568C;
        11'd1254   :   data <=16'h5681;
        11'd1255   :   data <=16'h5675;
        11'd1256   :   data <=16'h5669;
        11'd1257   :   data <=16'h565E;
        11'd1258   :   data <=16'h5652;
        11'd1259   :   data <=16'h5646;
        11'd1260   :   data <=16'h563B;

        11'd1261   :   data <=16'h562F;
        11'd1262   :   data <=16'h5624;
        11'd1263   :   data <=16'h5618;
        11'd1264   :   data <=16'h560C;
        11'd1265   :   data <=16'h5601;
        11'd1266   :   data <=16'h55F5;
        11'd1267   :   data <=16'h55EA;
        11'd1268   :   data <=16'h55DE;
        11'd1269   :   data <=16'h55D3;
        11'd1270   :   data <=16'h55C7;

        11'd1271   :   data <=16'h55BC;
        11'd1272   :   data <=16'h55B0;
        11'd1273   :   data <=16'h55A5;
        11'd1274   :   data <=16'h5599;
        11'd1275   :   data <=16'h558E;
        11'd1276   :   data <=16'h5582;
        11'd1277   :   data <=16'h5577;
        11'd1278   :   data <=16'h556C;
        11'd1279   :   data <=16'h5560;
        11'd1280   :   data <=16'h5555;

        default  :   data <= 16'h0000;
    endcase

endmodule
